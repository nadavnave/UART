`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:00:53 01/12/2021 
// Design Name: 
// Module Name:    UART_RX 
//	
//
//
//////////////////////////////////////////////////////////////////////////////////
module UART_RX(
    input serial_in,
    input x16_BAUD,
    input reset,
    output reg [7:0] Do,
    output reg valid,
    output reg error
    );


endmodule
